module BCDtoDecimal_300 (
    input clk,
    input reset,
    input [1199:0] bcd,
    output reg [3:0] dec
);

reg [8:0] index;
reg [3:0] temp_bcd;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        dec <= 4'd0;
        index <= 0;
    end 
    else if (index < 300) begin
        temp_bcd = bcd[(index * 4) +: 4];
        
        if (temp_bcd <= 4'd9) 
            dec <= temp_bcd;
        else
            dec <= 4'd0;

        index <= index + 1;
    end
end

endmodule
